`timescale 1ns / 1ps

module SerialSequenceDetector(
    input si,
    inout clk,
    output detected
    );


endmodule
